`timescale 1ns/1ps

module INSTRUCTION_FETCH(
	clk,
	rst,
	branch,
	branch_PC,
	//MEM_RW,
	
	PC,
	IR
);

input clk, rst;
input [31:0]branch_PC;
input [2:0] branch;
output reg 	[31:0] PC, IR;

//instruction memory
reg [31:0] instruction [300:0];

initial
begin
		instruction[ 0] = 32'b100011_00000_01000_00000_00000_000000;//lw $8,0($0)
		instruction[ 1] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 2] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 3] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 4] = 32'b000000_01000_00000_00011_00000_100000;	//add $3,$8,$2
		instruction[ 5] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 6] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 7] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 8] = 32'b000000_00011_00001_00011_00000_100000;//add $3,$3,$1
		instruction[ 9] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 10] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 11] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 12] = 32'b000000_00000_00001_00100_00000_100000;	//add $4,$0,$1
		instruction[ 13] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 14] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 15] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 16] = 32'b000000_00011_00010_00101_00000_100011;//4  div $5,$3,$2
		instruction[ 17] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 18] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 19] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 20] = 32'b000000_00100_00001_00100_00000_100000;//5  add $4,$4,$1
		instruction[ 21] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 22] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 23] = 32'b000000_00000_00000_00000_00000_100000;//
		//not yet
		instruction[ 24] = 32'b000100_00101_00100_00000_00000_001111;//6  beq $5,$4,15(to 40)
		instruction[ 25] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 26] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 27] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 28] = 32'b000000_00011_00100_00111_00000_100001;//7  mod $7,$3,$4
		instruction[ 29] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 30] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 31] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 32] = 32'b000100_00111_00000_11111_11111_100111;//8  beq $7,$0 -25(to 8)
		instruction[ 33] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 34] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 35] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 36] = 32'b000010_00000_00000_00000_00000_010100;//9 jump 20
		instruction[ 37] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 38] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 39] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 40] = 32'b101011_00000_00011_00000_00000_000001;//15 sw $3,1($0)
		instruction[ 41] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 42] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 43] = 32'b000000_00000_00000_00000_00000_100000;//
		
		///////////////////////////////////////////////////////////////////
		
		instruction[ 44] = 32'b100011_00000_01000_00000_00000_000000;//lw $8,0($0)
		instruction[ 45] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 46] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 47] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 48] = 32'b000000_01000_00000_00011_00000_100000;	//add $3,$8,$2
		instruction[ 49] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 50] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 51] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 52] = 32'b000000_00011_00001_00011_00000_100010;//add $3,$3,$1
		instruction[ 53] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 54] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 55] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 56] = 32'b000000_00000_00001_00100_00000_100000;	//add $4,$0,$1
		instruction[ 57] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 58] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 59] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 60] = 32'b000000_00011_00010_00101_00000_100011;//4  div $5,$3,$2
		instruction[ 61] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 62] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 63] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 64] = 32'b000000_00100_00001_00100_00000_100000;//5  add $4,$4,$1
		instruction[ 65] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 66] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 67] = 32'b000000_00000_00000_00000_00000_100000;//
		//not yet
		instruction[ 68] = 32'b000100_00101_00100_00000_00000_001111;//6  beq $5,$4,15(to 84)
		instruction[ 69] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 70] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 71] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 72] = 32'b000000_00011_00100_00111_00000_100001;//7  mod $7,$3,$4
		instruction[ 73] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 74] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 75] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 76] = 32'b000100_00111_00000_11111_11111_100111;//8  beq $7,$0 -25(to 52)
		instruction[ 77] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 78] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 79] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 80] = 32'b000010_00000_00000_00000_00001_000000;//9 jump 64
		instruction[ 81] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 82] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 83] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 84] = 32'b101011_00000_00011_00000_00000_000010;//15 sw $3,1($0)
		instruction[ 85] = 32'b000000_00000_00000_00000_00000_100000;	//
		instruction[ 86] = 32'b000000_00000_00000_00000_00000_100000;//
		instruction[ 87] = 32'b000000_00000_00000_00000_00000_100000;//
		
		instruction[ 88] = 32'b000010_00000_00000_00000_00001_011000;//9 jump 64
        instruction[ 89] = 32'b000000_00000_00000_00000_00000_100000;    //
        instruction[ 90] = 32'b000000_00000_00000_00000_00000_100000;//
        instruction[ 91] = 32'b000000_00000_00000_00000_00000_100000;//

end

//output instruction
always @(posedge clk or posedge rst)
begin
	if(rst)
		IR <= 32'd0;
	else
		IR <= instruction[PC[10:2]];
end

// output program counter
always @(posedge clk or posedge rst)
begin
	if(rst)
		PC <= 32'd0;
	else if(branch)
		PC <=branch_PC;
	else//add new PC address here, ex: branch, jump...
		PC <= PC+4;
end

endmodule